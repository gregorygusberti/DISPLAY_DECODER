LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DISPLAY_DECODER IS
	GENERIC (
		CAT: STD_LOGIC := '0'
	);
	PORT (
		DATA:  IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLANK: IN STD_LOGIC;
		TEST:  IN STD_LOGIC;
		
		--  A, B, C, D ...
		SEGM: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END DISPLAY_DECODER;

ARCHITECTURE ARCH OF DISPLAY_DECODER IS
	SIGNAL DC_O:     STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL PRE_OUT:  STD_LOGIC_VECTOR(6 DOWNTO 0);
	
	BEGIN
	
		SEGM <= PRE_OUT WHEN (CAT = '1') ELSE (NOT PRE_OUT);
	
		PRE_OUT <= "0000000" WHEN (BLANK = '1') ELSE "1111111" WHEN (TEST = '1') ELSE DC_O;
		
		WITH DATA SELECT
			DC_O <= "1111110" WHEN "0000",
					  "0110000" WHEN "0001",
					  "1101101" WHEN "0010",
					  "1111001" WHEN "0011",
					  "0110011" WHEN "0100",
					  "1011011" WHEN "0101",
					  "0011111" WHEN "0110",
					  "1110000" WHEN "0111",
					  "1111111" WHEN "1000",
					  "1110011" WHEN "1001",
					  "1001111" WHEN OTHERS;
					  
END ARCH;
					  
		